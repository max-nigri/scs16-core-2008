    0 => "00000000000000000000000000000000", 
    1 => "01101000000000000000000000000100", 
    2 => "01101000000000000000000001011001", 
    3 => "01101000000000000000000001011010", 
    4 => "00111000000100000000111111111111", 
    5 => "00111000000100110000000001000000", 
    6 => "00111000000100111000000001000001", 
    7 => "00011000000110001000000100001111", 
    8 => "00011000000110001000000000001111", 
    9 => "00011000000111010000000100001111", 
   10 => "00011000000111010000000000001111", 
   11 => "00011000000110011000000100000110", 
   12 => "00011000000110011000000000000111", 
   13 => "00011000000111100000000100000110", 
   14 => "00011000000111100000000000000111", 
   15 => "00111000000100110000000001000010", 
   16 => "00111000000100111000000001000011", 
   17 => "00111000000000001011000001100100", 
   18 => "00111000000010001011000100011110", 
   19 => "00111000000010010011000000011110", 
   20 => "00111000000100110000000001000110", 
   21 => "00111000000100111000000001001010", 
   22 => "00011100000111010000000100001111", 
   23 => "00011100000111010000000000001111", 
   24 => "00011100000110001000000100001111", 
   25 => "00011100000110001000000000001111", 
   26 => "00011100000111100000000100000110", 
   27 => "00011100000111100000000000000111", 
   28 => "00011100000110011000000100000110", 
   29 => "00011100000110011000000000000111", 
   30 => "00111000000100110000000001000010", 
   31 => "00111000000100111000000001000011", 
   32 => "00111100000000001011000001100100", 
   33 => "00111100000010001011000100011110", 
   34 => "00111100000010010011000000011110", 
   35 => "00111000000100110000000001000100", 
   36 => "00111000000100111000000001000101", 
   37 => "00111100001000001011000100011110", 
   38 => "00111100001000010011000000011110", 
   39 => "00111000000100010000000001011010", 
   40 => "00111000000100110000000000010100", 
   41 => "00111000000100111000000000011000", 
   42 => "01111000000100000000111110010000", 
   43 => "01111000000100000000111010010000", 
   44 => "00100000000110000010011100001111", 
   45 => "00100000000110000010011000001111", 
   46 => "00100000000111000010011100001111", 
   47 => "00100000000111000010011000001111", 
   48 => "00111000000100110000000000011110", 
   49 => "00111000000100111000000000100010", 
   50 => "00100000000110000010011100000110", 
   51 => "00100000000110000010011000000111", 
   52 => "00100000000111000010011100000110", 
   53 => "00100000000111000010011000000111", 
   54 => "01111000000000000010011000011110", 
   55 => "01111000000010000010011100011110", 
   56 => "01111000000010000010011000011110", 
   57 => "00111000000100010000000001011010", 
   58 => "00111000000100110000000000010100", 
   59 => "00111000000100111000000000011000", 
   60 => "01111100000100000000111110010000", 
   61 => "01111100000100000000111010010000", 
   62 => "00100100000110000010011100001111", 
   63 => "00100100000110000010011000001111", 
   64 => "00100100000111000010011100001111", 
   65 => "00100100000111000010011000001111", 
   66 => "00111000000100110000000000011110", 
   67 => "00111000000100111000000000100010", 
   68 => "00100100000110000010011100000110", 
   69 => "00100100000110000010011000000111", 
   70 => "00100100000111000010011100000110", 
   71 => "00100100000111000010011000000111", 
   72 => "01111100000000000010011000011110", 
   73 => "01111100000010000010011100011110", 
   74 => "01111100000010000010011000011110", 
   75 => "00111000000100110000000000110000", 
   76 => "00111000000100111000000000110100", 
   77 => "01111100001000000010011100011110", 
   78 => "01111100001000000010011000011110", 
   79 => "00111000000110011000000000110011", 
   80 => "00111000000100001000000001111111", 
   81 => "01010000000011111001011000000000", 
   82 => "10000000000111011110000001010101", 
   83 => "01011000000000000000000000000010", 
   84 => "01101000000000000000000001010110", 
   85 => "01011000000000000000000000000011", 
   86 => "00111000000100101000000000001010", 
   87 => "01101000000100000000000001011011", 
   88 => "10000000000111001111000001011000", 
   89 => "01110000000100000000000000000000", 
   90 => "01101000000000000000000000000100", 
   91 => "01001000000101001000010000000000", 
   92 => "00000000000000000000000000000000", 
   93 => "01110000000000000000000000000000", 
