    0 => "00000000000000000000000000000000", 
    1 => "01101000000000000000000000000100", 
    2 => "01101000000000000000000000001100", 
    3 => "01101000000000000000000000001101", 
    4 => "00111000000100000000111111111111", 
    5 => "01111000000000111000011011110000", 
    6 => "00111000000100110000000000010100", 
    7 => "00100100000110000110011100001111", 
    8 => "00000000000000000000000000000000", 
    9 => "00011100000110101000000100001111", 
   10 => "01101000000100000000000000001110", 
   11 => "10000000000111001111000000001011", 
   12 => "01110000000100000000000000000000", 
   13 => "01101000000000000000000000000100", 
   14 => "01001000000101001000010000000000", 
   15 => "00000000000000000000000000000000", 
   16 => "01110000000000000000000000000000", 
