    0 => "00000000000000000000000000000000", 
    1 => "00111000000100110000000000010000", 
    2 => "01111000000101000000011100001001", 
    3 => "01111000000101000000011100001001", 
    4 => "01111000000101100011111110000000", 
    5 => "00111000000100101000000000010100", 
    6 => "01001000000101100010100000000000", 
    7 => "00111000000100110000000000010001", 
    8 => "00011000000111001000000100001111", 
    9 => "00011000000111000000000100001111", 
   10 => "10000000000000111111100000001101", 
   11 => "00000000000000000000000000000000", 
   12 => "01101000000000000000000000010001", 
   13 => "10001000000000111001100000000000", 
   14 => "00100000000110000100011000001111", 
   15 => "10001000000000100100100000000001", 
   16 => "10101000000100000000000000000000", 
   17 => "01111000000000000001011000010001", 
   18 => "01111000000000000000011000010010", 
   19 => "00111000000000001011000000010000", 
   20 => "01001000000101001001100000000000", 
   21 => "10000000000000111111000000011000", 
   22 => "00000000000000000000000000000000", 
   23 => "01101000000000000000000000011011", 
   24 => "10001000000000111001100000000000", 
   25 => "00011000000110100000000000001111", 
   26 => "10101000000000000000000000000000", 
   27 => "01111000000000000001011000010000", 
   28 => "01111000000000000000011000010010", 
   29 => "10000000000111001111000000011101", 
   30 => "00000000000000000000000000000000", 
