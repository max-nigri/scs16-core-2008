    0 => "00000000000000000000000000000000", 
    1 => "01101000000000000000000000000100", 
    2 => "01101000000000000000000001000111", 
    3 => "01101000000000000000000001001000", 
    4 => "00111000000100000000111111111111", 
    5 => "01111000000000111000011011110000", 
    6 => "00111000000100101000000000000101", 
    7 => "10000000000101111001000000001001", 
    8 => "00111000000100001000000000000001", 
    9 => "10000000000101110001000000001011", 
   10 => "00111000000100001000000000000010", 
   11 => "00111000000100001000000000011110", 
   12 => "10000000000111001000000000001110", 
   13 => "00111000000100001000000000000001", 
   14 => "10000000000111001100000000010000", 
   15 => "00111000000100001000000000000010", 
   16 => "00111000000100001000000000101000", 
   17 => "10000000000111001000000000010100", 
   18 => "00111000000100001000000000000111", 
   19 => "01101000000000000000000000010101", 
   20 => "00111000000100001000000000001000", 
   21 => "10000000000111001100000000011000", 
   22 => "00111000000100001000000000001001", 
   23 => "01101000000000000000000000011001", 
   24 => "00111000000100001000000000001010", 
   25 => "10000000000111001000000000100000", 
   26 => "10000000000111001000100000011110", 
   27 => "10000000000111001001000000011101", 
   28 => "00111000000100001000000000001011", 
   29 => "00111000000100001000000000001100", 
   30 => "00111000000100001000000000001101", 
   31 => "01101000000000000000000000100001", 
   32 => "00111000000100001000000000001110", 
   33 => "10000000000111001011000000100100", 
   34 => "00111000000100001000000000010100", 
   35 => "01101000000000000000000000101110", 
   36 => "10000000000111001011100000100111", 
   37 => "00111000000100001000000000010101", 
   38 => "01101000000000000000000000101110", 
   39 => "10000000000111001100000000101010", 
   40 => "00111000000100001000000000010110", 
   41 => "01101000000000000000000000101110", 
   42 => "10000000000111001100100000101101", 
   43 => "00111000000100001000000000010111", 
   44 => "01101000000000000000000000101110", 
   45 => "00111000000100001000000000011000", 
   46 => "00111000000100010000000000101000", 
   47 => "10001000000000111010011000101000", 
   48 => "10000000000111011110000000110011", 
   49 => "00111000000100001000000000011110", 
   50 => "01101000000000000000000000110100", 
   51 => "00111000000100001000000000011111", 
   52 => "00111000000100010000000000101000", 
   53 => "10001000000000111010011000101000", 
   54 => "10000000000111011110000000111000", 
   55 => "00111000000100001000000000011110", 
   56 => "00111000000100010000000000101000", 
   57 => "10001000000000111010011000101000", 
   58 => "10000000000111011110100000111101", 
   59 => "00111000000100001000000000011110", 
   60 => "01101000000000000000000001000010", 
   61 => "10000000000111011101100001000000", 
   62 => "00111000000100001000000000011111", 
   63 => "01101000000000000000000001000010", 
   64 => "10000000000111011110000001000010", 
   65 => "00111000000100001000000000011111", 
   66 => "00111000000100010000000000110010", 
   67 => "10000000000010110000000001000101", 
   68 => "00111000000100010000000000111100", 
   69 => "00111000000100010000000001000110", 
   70 => "10000000000111001111000001000110", 
   71 => "01110000000100000000000000000000", 
   72 => "01101000000000000000000000000100", 
   73 => "01001000000101001000010000000000", 
   74 => "00000000000000000000000000000000", 
   75 => "01110000000000000000000000000000", 
